`include "dataflow.v"
module logic_gates_tb(input wire and_gate,or_gate, )
